----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    04:23:13 12/14/2009 
-- Design Name: 
-- Module Name:    vend_mach - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity vend_mach is
    Port ( switch : in  STD_LOGIC_VECTOR (1 downto 0);
           res_g : in  STD_LOGIC;
           res_l : in  STD_LOGIC;
           go : in  STD_LOGIC;
           item_price : in  STD_LOGIC_VECTOR (7 downto 0);
           change : out  STD_LOGIC_VECTOR (7 downto 0);
           disp : out  STD_LOGIC);
end vend_mach;

architecture Behavioral of vend_mach is

--type func is ()
type product is(gum,tofee,chocolate,lollypop);
signal avail_prod:product;
type price is array(0 to 3) of std_logic_vector(5 downto 0);
signal item_price: price<=(20,10,5,22);
type coin_typ is(one,two,five);
signal coin :coin_typ;
signal sum,change:STD_LOGIC_VECTOR (7 downto 0);

type state is (ini,ps,w,add,s4,s5);
signal nxt_state,cur_state: state;

begin

seq_log:	process(clk)
begin 
	if(clk='1' and clk'event)then
		cur_state<=nxt_state;
	end if;
end process;

comb_log:process(x,cur_state)
begin 
	case cur_state is
		WHEN s0 =>
			if(x='0')then 
				nxt_state<=s0;
				z<='0';
			else if(x='1')then 
				nxt_state<=s1;
				z<='0';
			end if;
			end if;
		
		when s1 =>
			if(x='0')then
				nxt_state<=s2;
			else if(x='1')then
				nxt_state<=s1;
			end if;
			end if;
		when s2 =>
			if(x='0')then
				nxt_state<=s0;
			else if(x='1')then
				nxt_state<=s3;
			end if;
			end if;
		when s3 =>
			if(x='0')then
				nxt_state<=s2;
			else if(x='1')then
				nxt_state<=s4;
			end if;
			end if;
		when s4 =>
			if(x='0')then
				nxt_state<=s5;
			else if(x='1')then
				nxt_state<=s1;
			end if;
			end if;
			
			when s5 =>
			
			nxt_state<=s0;
			if(x='1')then
			z<='1';
			end if;
			

		end case;
	end process;


end Behavioral;

